module adda(
			input			 ad_clk,
			input			 da_clk,
			input	[11:0]	 ad_data,
			output reg[11:0] da_data

);



endmodule